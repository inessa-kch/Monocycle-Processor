LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;



-----------------------------------------
ENTITY tb_Unite_de_Traitement IS
    ---------------------------------------

END ENTITY tb_Unite_de_Traitement;


